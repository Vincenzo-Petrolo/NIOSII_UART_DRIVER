-- niosii_system_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity niosii_system_tb is
end entity niosii_system_tb;

architecture rtl of niosii_system_tb is
	component niosii_system is
		port (
			clk_clk           : in  std_logic := 'X'; -- clk
			debug_pin_export  : out std_logic;        -- export
			pins_input_export : in  std_logic := 'X'; -- export
			reset_reset_n     : in  std_logic := 'X'  -- reset_n
		);
	end component niosii_system;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			sig_export : in std_logic_vector(0 downto 0) := (others => 'X')  -- export
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			sig_export : out std_logic_vector(0 downto 0)   -- export
		);
	end component altera_conduit_bfm_0002;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal niosii_system_inst_clk_bfm_clk_clk               : std_logic;                    -- niosii_system_inst_clk_bfm:clk -> [niosii_system_inst:clk_clk, niosii_system_inst_reset_bfm:clk]
	signal niosii_system_inst_debug_pin_export              : std_logic;                    -- niosii_system_inst:debug_pin_export -> niosii_system_inst_debug_pin_bfm:sig_export
	signal niosii_system_inst_pins_input_bfm_conduit_export : std_logic_vector(0 downto 0); -- niosii_system_inst_pins_input_bfm:sig_export -> niosii_system_inst:pins_input_export
	signal niosii_system_inst_reset_bfm_reset_reset         : std_logic;                    -- niosii_system_inst_reset_bfm:reset -> niosii_system_inst:reset_reset_n

begin
uart_tx : process
constant bit_time : TIME := 17us;
begin
niosii_system_inst_pins_input_bfm_conduit_export <= "1";
WAIT FOR 2ms; -- wait some time and send char 'U' corresponding to 0x55
niosii_system_inst_pins_input_bfm_conduit_export <= "0"; --glitch
WAIT FOR 5us;
niosii_system_inst_pins_input_bfm_conduit_export <= "1";
WAIT FOR 40us;
niosii_system_inst_pins_input_bfm_conduit_export <= "0";--start bit
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "1"; --lsb
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "0";
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "1";
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "0";
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "1";
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "0";
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "1";
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "0";--msb
WAIT FOR bit_time;
niosii_system_inst_pins_input_bfm_conduit_export <= "1"; --STOP
end process;
	niosii_system_inst : component niosii_system
		port map (
			clk_clk           => niosii_system_inst_clk_bfm_clk_clk,                  --        clk.clk
			debug_pin_export  => niosii_system_inst_debug_pin_export,                 --  debug_pin.export
			pins_input_export => niosii_system_inst_pins_input_bfm_conduit_export(0), -- pins_input.export
			reset_reset_n     => niosii_system_inst_reset_bfm_reset_reset             --      reset.reset_n
		);

	niosii_system_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 100000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => niosii_system_inst_clk_bfm_clk_clk  -- clk.clk
		);

--	niosii_system_inst_debug_pin_bfm : component altera_conduit_bfm
--		port map (
--			sig_export(0) => niosii_system_inst_debug_pin_export  -- conduit.export
--		);
--
--	niosii_system_inst_pins_input_bfm : component altera_conduit_bfm_0002
--		port map (
--			sig_export => niosii_system_inst_pins_input_bfm_conduit_export  -- conduit.export
--		);

	niosii_system_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => niosii_system_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => niosii_system_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of niosii_system_tb
